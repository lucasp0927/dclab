module rsa (/*AUTOARG*/
	    // Outputs
	    ready, data_o,
	    // Inputs
	    clk, reset, we, oe, start, reg_sel, addr, data_i
	    );
   input clk,reset,we,oe,start;
   input [1:0] reg_sel;
   input [4:0] addr;
   input [7:0] data_i;
   output      ready;
   output [7:0] data_o;
   integer 	addr_num;
   reg [255:0] 	a[3:0]; //a[0] = a[1]^a[2] mod a[3]
   /*AUTOREG*/
   // Beginning of automatic regs (for this module's undeclared outputs)
   reg [7:0] 	data_o;
   reg 		ready;
   // End of automatics
   /*AUTOWIRE*/

   ////////////////////////////////////////////////////////////////////////////////////////////////////
   //    io
   ////////////////////////////////////////////////////////////////////////////////////////////////////
   always @(posedge clk) begin
      if ((we==0) || (oe==0)) begin
	 case (reg_sel)
	   2'd0:
	     begin
		case (addr)
		  5'd0: a[0][1*8-1:0]<=data_i;
		  5'd1: a[0][2*8-1:1*8]<=data_i;
		  5'd2: a[0][3*8-1:2*8]<=data_i;
		  5'd3: a[0][4*8-1:3*8]<=data_i;
		  5'd4: a[0][5*8-1:4*8]<=data_i;
		  5'd5: a[0][6*8-1:5*8]<=data_i;
		  5'd6: a[0][7*8-1:6*8]<=data_i;
		  5'd7: a[0][8*8-1:7*8]<=data_i;
		  5'd8: a[0][9*8-1:8*8]<=data_i;
		  5'd9: a[0][10*8-1:9*8]<=data_i;
		  5'd10: a[0][11*8-1:10*8]<=data_i;
		  5'd11: a[0][12*8-1:11*8]<=data_i;
		  5'd12: a[0][13*8-1:12*8]<=data_i;
		  5'd13: a[0][14*8-1:13*8]<=data_i;
		  5'd14: a[0][15*8-1:14*8]<=data_i;
		  5'd15: a[0][16*8-1:15*8]<=data_i;
		  5'd16: a[0][17*8-1:16*8]<=data_i;
		  5'd17: a[0][18*8-1:17*8]<=data_i;
		  5'd18: a[0][19*8-1:18*8]<=data_i;
		  5'd19: a[0][20*8-1:19*8]<=data_i;
		  5'd20: a[0][21*8-1:20*8]<=data_i;
		  5'd21: a[0][22*8-1:21*8]<=data_i;
		  5'd22: a[0][23*8-1:22*8]<=data_i;
		  5'd23: a[0][24*8-1:23*8]<=data_i;
		  5'd24: a[0][25*8-1:24*8]<=data_i;
		  5'd25: a[0][26*8-1:25*8]<=data_i;
		  5'd26: a[0][27*8-1:26*8]<=data_i;
		  5'd27: a[0][28*8-1:27*8]<=data_i;
		  5'd28: a[0][29*8-1:28*8]<=data_i;
		  5'd29: a[0][30*8-1:29*8]<=data_i;
		  5'd30: a[0][31*8-1:30*8]<=data_i;
		  5'd31: a[0][32*8-1:31*8]<=data_i;
		endcase
	     end
	   2'd1:
	     begin
		case (addr)
		  5'd0: a[1][1*8-1:0]<=data_i;
		  5'd1: a[1][2*8-1:1*8]<=data_i;
		  5'd2: a[1][3*8-1:2*8]<=data_i;
		  5'd3: a[1][4*8-1:3*8]<=data_i;
		  5'd4: a[1][5*8-1:4*8]<=data_i;
		  5'd5: a[1][6*8-1:5*8]<=data_i;
		  5'd6: a[1][7*8-1:6*8]<=data_i;
		  5'd7: a[1][8*8-1:7*8]<=data_i;
		  5'd8: a[1][9*8-1:8*8]<=data_i;
		  5'd9: a[1][10*8-1:9*8]<=data_i;
		  5'd10: a[1][11*8-1:10*8]<=data_i;
		  5'd11: a[1][12*8-1:11*8]<=data_i;
		  5'd12: a[1][13*8-1:12*8]<=data_i;
		  5'd13: a[1][14*8-1:13*8]<=data_i;
		  5'd14: a[1][15*8-1:14*8]<=data_i;
		  5'd15: a[1][16*8-1:15*8]<=data_i;
		  5'd16: a[1][17*8-1:16*8]<=data_i;
		  5'd17: a[1][18*8-1:17*8]<=data_i;
		  5'd18: a[1][19*8-1:18*8]<=data_i;
		  5'd19: a[1][20*8-1:19*8]<=data_i;
		  5'd20: a[1][21*8-1:20*8]<=data_i;
		  5'd21: a[1][22*8-1:21*8]<=data_i;
		  5'd22: a[1][23*8-1:22*8]<=data_i;
		  5'd23: a[1][24*8-1:23*8]<=data_i;
		  5'd24: a[1][25*8-1:24*8]<=data_i;
		  5'd25: a[1][26*8-1:25*8]<=data_i;
		  5'd26: a[1][27*8-1:26*8]<=data_i;
		  5'd27: a[1][28*8-1:27*8]<=data_i;
		  5'd28: a[1][29*8-1:28*8]<=data_i;
		  5'd29: a[1][30*8-1:29*8]<=data_i;
		  5'd30: a[1][31*8-1:30*8]<=data_i;
		  5'd31: a[1][32*8-1:31*8]<=data_i;
		endcase
	     end
	   2'd2:
	     begin
		case (addr)
		  5'd0: a[2][1*8-1:0]<=data_i;
		  5'd1: a[2][2*8-1:1*8]<=data_i;
		  5'd2: a[2][3*8-1:2*8]<=data_i;
		  5'd3: a[2][4*8-1:3*8]<=data_i;
		  5'd4: a[2][5*8-1:4*8]<=data_i;
		  5'd5: a[2][6*8-1:5*8]<=data_i;
		  5'd6: a[2][7*8-1:6*8]<=data_i;
		  5'd7: a[2][8*8-1:7*8]<=data_i;
		  5'd8: a[2][9*8-1:8*8]<=data_i;
		  5'd9: a[2][10*8-1:9*8]<=data_i;
		  5'd10: a[2][11*8-1:10*8]<=data_i;
		  5'd11: a[2][12*8-1:11*8]<=data_i;
		  5'd12: a[2][13*8-1:12*8]<=data_i;
		  5'd13: a[2][14*8-1:13*8]<=data_i;
		  5'd14: a[2][15*8-1:14*8]<=data_i;
		  5'd15: a[2][16*8-1:15*8]<=data_i;
		  5'd16: a[2][17*8-1:16*8]<=data_i;
		  5'd17: a[2][18*8-1:17*8]<=data_i;
		  5'd18: a[2][19*8-1:18*8]<=data_i;
		  5'd19: a[2][20*8-1:19*8]<=data_i;
		  5'd20: a[2][21*8-1:20*8]<=data_i;
		  5'd21: a[2][22*8-1:21*8]<=data_i;
		  5'd22: a[2][23*8-1:22*8]<=data_i;
		  5'd23: a[2][24*8-1:23*8]<=data_i;
		  5'd24: a[2][25*8-1:24*8]<=data_i;
		  5'd25: a[2][26*8-1:25*8]<=data_i;
		  5'd26: a[2][27*8-1:26*8]<=data_i;
		  5'd27: a[2][28*8-1:27*8]<=data_i;
		  5'd28: a[2][29*8-1:28*8]<=data_i;
		  5'd29: a[2][30*8-1:29*8]<=data_i;
		  5'd30: a[2][31*8-1:30*8]<=data_i;
		  5'd31: a[2][32*8-1:31*8]<=data_i;
		endcase
	     end
	   2'd3:
	     begin
		;
		
	     end
	   default:
	     begin
		;
		
	     end
	 endcase // case (reg_sel)
      end
   end 

endmodule

