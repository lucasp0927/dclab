module io (/*AUTOARG*/
   // Outputs
   a,
   // Inputs
   addr, data_i
   );

   input [4:0] addr;
   input [7:0] data_i;
   output [255:0] a;
	 
endmodule
